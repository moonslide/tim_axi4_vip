`ifndef AXI4_TC_005_EXHAUSTIVE_RANDOM_READS_VIRTUAL_SEQ_INCLUDED_
`define AXI4_TC_005_EXHAUSTIVE_RANDOM_READS_VIRTUAL_SEQ_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: axi4_tc_005_exhaustive_random_reads_virtual_seq
// Test Case 5: Exhaustive Randomized Read & Boundary Verification
//--------------------------------------------------------------------------------------------
class axi4_tc_005_exhaustive_random_reads_virtual_seq extends axi4_virtual_base_seq;
  
  `uvm_object_utils(axi4_tc_005_exhaustive_random_reads_virtual_seq)

  // Random read sequences for each master
  axi4_master_bk_read_seq random_read_seq_h[10];
  
  // Slave sequences
  axi4_slave_bk_read_seq axi4_slave_read_seq_h[10];

  // Configuration parameters
  int NUM_TRANSACTIONS_PER_PAIR = 2; // Reduced for practical simulation time
  int total_transactions = 0;
  int boundary_crossings = 0;

  extern function new(string name = "axi4_tc_005_exhaustive_random_reads_virtual_seq");
  extern task body();
  extern task setup_slave_sequences();
  extern task execute_exhaustive_matrix_reads();
  extern task check_4k_boundary_crossing(bit [63:0] start_addr, int len, int size);

endclass : axi4_tc_005_exhaustive_random_reads_virtual_seq

function axi4_tc_005_exhaustive_random_reads_virtual_seq::new(string name = "axi4_tc_005_exhaustive_random_reads_virtual_seq");
  super.new(name);
endfunction : new

task axi4_tc_005_exhaustive_random_reads_virtual_seq::body();
  
  `uvm_info("TC005_VSEQ", "Starting TC005 Exhaustive Randomized Read Matrix Test", UVM_NONE);
  `uvm_info("TC005_VSEQ", $sformatf("Testing 10x10 Master-Slave Matrix (%0d transactions per pair)", NUM_TRANSACTIONS_PER_PAIR), UVM_NONE);
  
  super.body();
  
  // Create read sequence handles
  foreach(random_read_seq_h[i]) begin
    random_read_seq_h[i] = axi4_master_bk_read_seq::type_id::create($sformatf("random_read_seq_h[%0d]", i));
  end
  
  setup_slave_sequences();
  execute_exhaustive_matrix_reads();
  
  `uvm_info("TC005_VSEQ", "========================================", UVM_NONE);
  `uvm_info("TC005_VSEQ", "TC005 Exhaustive Random Read Matrix COMPLETE", UVM_NONE);
  `uvm_info("TC005_VSEQ", $sformatf("Total transactions: %0d", total_transactions), UVM_NONE);
  `uvm_info("TC005_VSEQ", $sformatf("4K boundary crossings detected: %0d", boundary_crossings), UVM_NONE);
  `uvm_info("TC005_VSEQ", "========================================", UVM_NONE);
  
endtask : body

task axi4_tc_005_exhaustive_random_reads_virtual_seq::setup_slave_sequences();
  
  foreach(axi4_slave_read_seq_h[i]) begin
    axi4_slave_read_seq_h[i] = axi4_slave_bk_read_seq::type_id::create($sformatf("axi4_slave_read_seq_h[%0d]", i));
  end
  
  // Start slave sequences for all 10 slaves with timeout protection (reduced repeat counts)
  fork
    begin : SLAVE_RESPONSES
      fork
        begin : SLAVE_S0_HANDLER
          repeat(10) axi4_slave_read_seq_h[0].start(p_sequencer.axi4_slave_read_seqr_h_all[0]); // S0
        end
        begin : SLAVE_S1_HANDLER  
          repeat(10) axi4_slave_read_seq_h[1].start(p_sequencer.axi4_slave_read_seqr_h_all[1]); // S1
        end
        begin : SLAVE_S2_HANDLER
          repeat(10) axi4_slave_read_seq_h[2].start(p_sequencer.axi4_slave_read_seqr_h_all[2]); // S2
        end
        begin : SLAVE_S3_HANDLER
          repeat(10) axi4_slave_read_seq_h[3].start(p_sequencer.axi4_slave_read_seqr_h_all[3]); // S3
        end
        begin : SLAVE_S4_HANDLER
          repeat(10) axi4_slave_read_seq_h[4].start(p_sequencer.axi4_slave_read_seqr_h_all[4]); // S4
        end
        begin : SLAVE_S5_HANDLER
          repeat(10) axi4_slave_read_seq_h[5].start(p_sequencer.axi4_slave_read_seqr_h_all[5]); // S5
        end
        begin : SLAVE_S6_HANDLER
          repeat(10) axi4_slave_read_seq_h[6].start(p_sequencer.axi4_slave_read_seqr_h_all[6]); // S6
        end
        begin : SLAVE_S7_HANDLER
          repeat(10) axi4_slave_read_seq_h[7].start(p_sequencer.axi4_slave_read_seqr_h_all[7]); // S7
        end
        begin : SLAVE_S8_HANDLER
          repeat(10) axi4_slave_read_seq_h[8].start(p_sequencer.axi4_slave_read_seqr_h_all[8]); // S8
        end
        begin : SLAVE_S9_HANDLER
          repeat(10) axi4_slave_read_seq_h[9].start(p_sequencer.axi4_slave_read_seqr_h_all[9]); // S9
        end
        begin : SLAVE_TIMEOUT
          #25000; // 25000 time units timeout for slave sequences
          `uvm_info("TC005_VSEQ", "Slave sequence timeout reached - ending slave responses", UVM_MEDIUM);
        end
      join_any
    end
  join_none
  
endtask : setup_slave_sequences

task axi4_tc_005_exhaustive_random_reads_virtual_seq::execute_exhaustive_matrix_reads();
  
  string expected_resp; // Declare string variable outside the loops
  
  `uvm_info("TC005_VSEQ", "Executing exhaustive 10x10 Master-Slave read matrix", UVM_MEDIUM);
  
  // Test every master-slave pairing (10x10 = 100 combinations)
  for (int master_id = 0; master_id < 10; master_id++) begin
    for (int slave_id = 0; slave_id < 10; slave_id++) begin
      
      `uvm_info("TC005_VSEQ", 
        $sformatf("Testing M%0d → S%0d pairing (%0d transactions)", 
        master_id, slave_id, NUM_TRANSACTIONS_PER_PAIR), UVM_MEDIUM);
      
      // Execute multiple random read transactions for this master-slave pair
      for (int trans = 0; trans < NUM_TRANSACTIONS_PER_PAIR; trans++) begin
        
        axi4_master_tx req;
        bit [63:0] slave_base_addr;
        bit [63:0] slave_end_addr;
        
        // Define slave address ranges based on claude.md
        case(slave_id)
          0: begin slave_base_addr = 64'h1000_0000; slave_end_addr = 64'h1FFF_FFFF; end // S0: DDR Secure Kernel
          1: begin slave_base_addr = 64'h2000_0000; slave_end_addr = 64'h2FFF_FFFF; end // S1: DDR Non-Secure User
          2: begin slave_base_addr = 64'h3000_0000; slave_end_addr = 64'h3FFF_FFFF; end // S2: DDR Shared Buffer
          3: begin slave_base_addr = 64'h4000_0000; slave_end_addr = 64'h4FFF_FFFF; end // S3: Illegal Address Hole
          4: begin slave_base_addr = 64'h5000_0000; slave_end_addr = 64'h5FFF_FFFF; end // S4: XOM Instruction-Only
          5: begin slave_base_addr = 64'h6000_0000; slave_end_addr = 64'h6FFF_FFFF; end // S5: RO Peripheral
          6: begin slave_base_addr = 64'h7000_0000; slave_end_addr = 64'h7FFF_FFFF; end // S6: Privileged-Only
          7: begin slave_base_addr = 64'h8000_0000; slave_end_addr = 64'h8FFF_FFFF; end // S7: Secure-Only
          8: begin slave_base_addr = 64'h9000_0000; slave_end_addr = 64'h9FFF_FFFF; end // S8: Scratchpad
          9: begin slave_base_addr = 64'hA000_0000; slave_end_addr = 64'hAFFF_FFFF; end // S9: Attribute Monitor
          default: begin slave_base_addr = 64'h0; slave_end_addr = 64'hFFFF_FFFF; end
        endcase
        
        // Create and randomize transaction
        req = axi4_master_tx::type_id::create("req");
        
        if(!req.randomize() with {
          req.tx_type == READ;
          req.transfer_type == BLOCKING_READ;
          req.araddr >= slave_base_addr && req.araddr <= slave_end_addr;
          req.arsize inside {READ_1_BYTE, READ_2_BYTES, READ_4_BYTES, READ_8_BYTES};
          req.arlen inside {4'h0, 4'h1, 4'h3, 4'h7, 4'hF}; // Various burst lengths
          req.arburst == READ_INCR;
          
          // Master-specific AxPROT constraints (simplified)
          if (master_id == 0) req.arprot == 3'b000; // M0: Secure CPU
          else if (master_id == 1) req.arprot == 3'b111; // M1: Non-secure CPU
          else if (master_id == 2) req.arprot == 3'b100; // M2: Instruction fetch
          else req.arprot inside {3'b000, 3'b111, 3'b110}; // Other masters
          
        }) begin
          `uvm_fatal("TC005_VSEQ", $sformatf("Randomization failed for M%0d→S%0d transaction %0d", master_id, slave_id, trans));
        end
        
        // Check for 4K boundary crossings
        check_4k_boundary_crossing(req.araddr, req.arlen, req.arsize);
        
        // Generate expected response based on master-slave access matrix
        expected_resp = "VARY"; // Default - depends on access matrix
        case ({master_id, slave_id})
          {4'd0, 4'd0}: expected_resp = "OKAY";  // M0→S0: Secure CPU to secure region
          {4'd1, 4'd0}: expected_resp = "DECERR"; // M1→S0: Non-secure to secure region
          {4'd2, 4'd4}: expected_resp = "OKAY";  // M2→S4: Instruction fetch to XOM
          {4'd7, 4'd4}: expected_resp = "SLVERR"; // M7→S4: Data access to instruction-only
          // Add more specific cases based on claude.md matrix...
          default: expected_resp = "MATRIX"; // Check full access matrix
        endcase
        
        // Execute the transaction - create new sequence instance for each transaction
        fork
          begin
            axi4_master_bk_read_seq temp_read_seq;
            temp_read_seq = axi4_master_bk_read_seq::type_id::create($sformatf("temp_read_seq_m%0d_s%0d_t%0d", master_id, slave_id, trans));
            temp_read_seq.start(p_sequencer.axi4_master_read_seqr_h_all[master_id]);
            total_transactions++;
          end
        join_none
        
        if (trans % 10 == 0) begin
          `uvm_info("TC005_VSEQ", 
            $sformatf("M%0d→S%0d: %0d/%0d transactions (Expect: %s)", 
            master_id, slave_id, trans, NUM_TRANSACTIONS_PER_PAIR, expected_resp), UVM_DEBUG);
        end
        
        #1; // Small delay between transactions
      end
      
      `uvm_info("TC005_VSEQ", 
        $sformatf("Completed M%0d→S%0d pairing", master_id, slave_id), UVM_MEDIUM);
      
      #10; // Inter-pairing delay
    end
  end
  
  // Wait for all transactions to complete with timeout protection
  fork
    begin : WAIT_FOR_COMPLETION
      wait fork;
    end
    begin : COMPLETION_TIMEOUT
      #50000; // 50000 time units timeout for all transactions to complete
      `uvm_warning("TC005_VSEQ", "Transaction completion timeout reached - proceeding with test completion");
    end
  join_any
  
  // Disable timeout thread if operations completed first
  disable COMPLETION_TIMEOUT;
  
  #2000;
  
  `uvm_info("TC005_VSEQ", "Exhaustive matrix read test completed", UVM_MEDIUM);
  
endtask : execute_exhaustive_matrix_reads

task axi4_tc_005_exhaustive_random_reads_virtual_seq::check_4k_boundary_crossing(bit [63:0] start_addr, int len, int size);
  
  bit [63:0] end_addr;
  bit [63:0] start_4k_boundary;
  bit [63:0] end_4k_boundary;
  int bytes_per_beat;
  
  // Calculate bytes per beat based on size
  case(size)
    0: bytes_per_beat = 1;  // READ_1_BYTE
    1: bytes_per_beat = 2;  // READ_2_BYTES
    2: bytes_per_beat = 4;  // READ_4_BYTES
    3: bytes_per_beat = 8;  // READ_8_BYTES
    default: bytes_per_beat = 4;
  endcase
  
  // Calculate end address of burst
  end_addr = start_addr + ((len + 1) * bytes_per_beat) - 1;
  
  // Calculate 4K boundaries
  start_4k_boundary = start_addr >> 12; // Divide by 4096
  end_4k_boundary = end_addr >> 12;     // Divide by 4096
  
  // Check if burst crosses 4K boundary
  if (start_4k_boundary != end_4k_boundary) begin
    boundary_crossings++;
    `uvm_warning("TC005_4K_BOUNDARY", 
      $sformatf("4K boundary crossing detected: Start=0x%16h, End=0x%16h, Len=%0d, Size=%0d", 
      start_addr, end_addr, len, size));
  end
  
endtask : check_4k_boundary_crossing

`endif