`ifndef AXI4_EXCEPTION_CLK_RESET_TESTS_INCLUDED_
`define AXI4_EXCEPTION_CLK_RESET_TESTS_INCLUDED_

//=============================================================================================
// File: axi4_exception_clk_reset_tests.sv
// Description: Clock and Reset Exception Tests for AXI4 Protocol
//
// This file contains test cases that inject clock frequency changes and reset events
// during active AXI4 transfers to test system resilience and recovery capabilities.
//
// TEST CASES INCLUDED:
// 1. axi4_exception_clk_freq_change_test
//    - Changes clock frequency during active transfers
//    - Tests system behavior with varying clock speeds
//    - Verifies data integrity across frequency transitions
//    - Frequency scaling: 0.5x to 3.0x of nominal
//    - Number of changes: 1-10 events (random)
//
// 2. axi4_exception_reset_terminate_test
//    - Asserts reset during active transfers
//    - Tests proper transaction abandonment
//    - Verifies system recovery after reset
//    - Reset duration: 1-10 cycles (random)
//    - Number of resets: 1-8 events (random)
//
// 3. axi4_exception_clk_reset_combined_test
//    - Combines clock frequency changes with reset events
//    - Tests system under combined stress scenarios
//    - Verifies recovery from simultaneous exceptions
//    - Mixed events: 3-15 total (random)
//
// 4. axi4_exception_continuous_clk_change_test
//    - Continuously varies clock frequency throughout test
//    - Tests system stability under constant frequency variation
//    - Change probability: 5-30% per interval
//    - Test duration: 5-20 microseconds
//
// COMMON FEATURES:
// - Random timing of exception events
// - Recovery verification after each event
// - Protocol compliance checking during exceptions
// - Performance metrics collection
// - Support for all bus matrix modes: NONE (1x1), BASE (4x4), ENHANCED (10x10)
//
// EXCEPTION PARAMETERS:
// - Clock frequency factors: 0.5x, 0.75x, 1.0x, 1.25x, 1.5x, 2.0x, 3.0x
// - Reset phases: Address, Data, Response, or Idle
// - Recovery timeout: Configurable (default 100 cycles)
// - Deadlock/livelock detection during exceptions
//
// USAGE IN REGRESSION:
// These tests are included in both error_inject.list and axi4_transfers_regression.list
// with run_cnt=3-5 for each bus matrix mode to ensure thorough exception coverage.
//=============================================================================================

//--------------------------------------------------------------------------------------------
// Class: axi4_exception_clk_freq_change_test
// Description:
// This test performs multiple clock frequency changes during active transfers.
// - Number of changes: 1-10 events (random)
// - Frequency scaling: 0.5x to 3.0x (random)
// - Change timing: During transfer or idle (random)
// - Hold duration: 5-100 cycles per frequency (random)
// - Recovery testing: Verifies proper recovery after frequency changes
// - Supports all bus matrix modes (NONE/1x1, BASE/4x4, ENHANCED/10x10)
//--------------------------------------------------------------------------------------------
class axi4_exception_clk_freq_change_test extends axi4_error_inject_base_test;
  `uvm_component_utils(axi4_exception_clk_freq_change_test)

  extern function new(string name = "axi4_exception_clk_freq_change_test", uvm_component parent = null);
  extern function void build_phase(uvm_phase phase);
  extern virtual function void setup_axi4_env_cfg();
  extern task run_phase(uvm_phase phase);
  extern function void report_phase(uvm_phase phase);

endclass : axi4_exception_clk_freq_change_test

function axi4_exception_clk_freq_change_test::new(string name = "axi4_exception_clk_freq_change_test", uvm_component parent = null);
  super.new(name, parent);
endfunction : new

function void axi4_exception_clk_freq_change_test::build_phase(uvm_phase phase);
  super.build_phase(phase);
  
  // Configure test for clock frequency exceptions
  uvm_config_db#(bit)::set(this, "*", "enable_exceptions", 1);
  uvm_config_db#(bit)::set(this, "*", "clk_freq_exception", 1);
  uvm_config_db#(bit)::set(this, "*", "randomize_freq_change", 1);
  uvm_config_db#(int)::set(this, "*", "max_freq_changes", 10);
  
  `uvm_info(get_type_name(), "Build phase completed for Clock Frequency Change Exception test", UVM_LOW)
endfunction : build_phase

function void axi4_exception_clk_freq_change_test::setup_axi4_env_cfg();
  // Call parent implementation first
  super.setup_axi4_env_cfg();
  
  // Enable frequency checker for this test
  axi4_env_cfg_h.has_freq_checker = 1;
  
  // Configure expected frequency changes for the checker
  // The test performs 1-10 random frequency changes
  uvm_config_db#(int)::set(this, "*", "expected_freq_changes", 10);
  
  `uvm_info(get_type_name(), "Enabled frequency checker for clock frequency change test", UVM_MEDIUM)
endfunction : setup_axi4_env_cfg

task axi4_exception_clk_freq_change_test::run_phase(uvm_phase phase);
  axi4_master_exception_clk_freq_seq clk_freq_seq[];
  int active_masters;
  int num_freq_events = 5;
  
  phase.raise_objection(this);
  
  // Determine active masters based on bus matrix mode
  case(test_config.bus_matrix_mode)
    axi4_bus_matrix_ref::NONE: active_masters = 1;
    axi4_bus_matrix_ref::BASE_BUS_MATRIX: active_masters = 4;
    axi4_bus_matrix_ref::BUS_ENHANCED_MATRIX: active_masters = test_config.num_masters;
  endcase
  
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  `uvm_info(get_type_name(), "Starting Clock Frequency Change Exception Test", UVM_LOW)
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  `uvm_info(get_type_name(), "Test Description:", UVM_LOW)
  `uvm_info(get_type_name(), "  - Multiple frequency changes (1-10 events)", UVM_LOW)
  `uvm_info(get_type_name(), "  - Frequency scaling: 0.5x to 3.0x", UVM_LOW)
  `uvm_info(get_type_name(), "  - Random timing during transfers", UVM_LOW)
  `uvm_info(get_type_name(), "  - Tests sampling error detection", UVM_LOW)
  `uvm_info(get_type_name(), $sformatf("  - Bus Matrix Mode: %s with %0dx%0d configuration", 
            test_config.bus_matrix_mode.name(), test_config.num_masters, test_config.num_slaves), UVM_LOW)
  `uvm_info(get_type_name(), $sformatf("  - Testing %0d active masters", active_masters), UVM_LOW)
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  
  // Configure expected frequency changes for the checker
  if(axi4_env_h.axi4_freq_checker_h != null) begin
    // Don't set strict expectations, just monitor
    axi4_env_h.axi4_freq_checker_h.expected_freq_changes = 0;  // 0 means no strict checking
  end
  
  // Create sequences for each active master
  clk_freq_seq = new[active_masters];
  
  // Run frequency change sequences on multiple masters
  fork
    begin
      for(int m = 0; m < active_masters; m++) begin
        automatic int master_id = m;
        fork
          begin
            clk_freq_seq[master_id] = axi4_master_exception_clk_freq_seq::type_id::create($sformatf("clk_freq_seq_%0d", master_id));
            
            // Randomize for this master
            if(!clk_freq_seq[master_id].randomize() with {
              num_freq_changes inside {[1:3]};
            }) begin
              `uvm_error(get_type_name(), $sformatf("Failed to randomize freq sequence for master %0d", master_id))
            end
            
            // Add some delay to stagger the frequency changes
            #(master_id * 100ns);
            
            `uvm_info(get_type_name(), $sformatf("Starting freq changes on master %0d", master_id), UVM_LOW)
            
            if (test_config.num_masters > master_id) begin
              clk_freq_seq[master_id].start(axi4_env_h.axi4_virtual_seqr_h.axi4_master_write_seqr_h_all[master_id]);
            end
          end
        join_none
      end
      
      // Wait for all masters to complete
      wait fork;
    end
  join
  
  // Wait for completion
  #1000ns;
  
  phase.drop_objection(this);
  
endtask : run_phase

function void axi4_exception_clk_freq_change_test::report_phase(uvm_phase phase);
  uvm_report_server svr;
  super.report_phase(phase);
  
  svr = uvm_report_server::get_server();
  
  if(svr.get_severity_count(UVM_FATAL) + svr.get_severity_count(UVM_ERROR) == 0) begin
    `uvm_info(get_type_name(), "===============================================", UVM_LOW)
    `uvm_info(get_type_name(), "Clock Frequency Change Exception Test PASSED", UVM_LOW)
    `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  end else begin
    `uvm_info(get_type_name(), "===============================================", UVM_LOW)
    `uvm_info(get_type_name(), "Clock Frequency Change Exception Test FAILED", UVM_LOW)
    `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  end
endfunction : report_phase

//--------------------------------------------------------------------------------------------
// Class: axi4_exception_reset_terminate_test
// Description:
// This test performs reset assertion during active transfers.
// - Number of resets: 1-8 events (random)
// - Reset duration: 1-10 cycles (random)
// - Reset phases: Address, Data, Response, or Idle (random)
// - Transfer abandonment: Verifies proper cleanup
// - Recovery testing: Ensures system recovers after reset
// - Supports all bus matrix modes (NONE/1x1, BASE/4x4, ENHANCED/10x10)
//--------------------------------------------------------------------------------------------
class axi4_exception_reset_terminate_test extends axi4_error_inject_base_test;
  `uvm_component_utils(axi4_exception_reset_terminate_test)

  extern function new(string name = "axi4_exception_reset_terminate_test", uvm_component parent = null);
  extern function void build_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);

endclass : axi4_exception_reset_terminate_test

function axi4_exception_reset_terminate_test::new(string name = "axi4_exception_reset_terminate_test", uvm_component parent = null);
  super.new(name, parent);
endfunction : new

function void axi4_exception_reset_terminate_test::build_phase(uvm_phase phase);
  super.build_phase(phase);
  
  // Configure test for reset termination exceptions
  uvm_config_db#(bit)::set(this, "*", "enable_exceptions", 1);
  uvm_config_db#(bit)::set(this, "*", "reset_terminate", 1);
  uvm_config_db#(bit)::set(this, "*", "verify_abandonment", 1);
  uvm_config_db#(int)::set(this, "*", "max_reset_events", 8);
  
  `uvm_info(get_type_name(), "Build phase completed for Reset Terminate test", UVM_LOW)
endfunction : build_phase

task axi4_exception_reset_terminate_test::run_phase(uvm_phase phase);
  axi4_master_exception_reset_terminate_seq reset_seq;
  
  phase.raise_objection(this);
  
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  `uvm_info(get_type_name(), "Starting Reset Termination Exception Test", UVM_LOW)
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  `uvm_info(get_type_name(), "Test Description:", UVM_LOW)
  `uvm_info(get_type_name(), "  - Multiple reset events (1-8 times)", UVM_LOW)
  `uvm_info(get_type_name(), "  - Reset during different phases", UVM_LOW)
  `uvm_info(get_type_name(), "  - Verifies transfer abandonment", UVM_LOW)
  `uvm_info(get_type_name(), "  - Tests recovery after reset", UVM_LOW)
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  
  // Run the reset termination sequence on first master
  reset_seq = axi4_master_exception_reset_terminate_seq::type_id::create("reset_seq");
  
  // Randomize to get multiple reset events (3-5 events for testing)
  if(!reset_seq.randomize() with {
    num_reset_events inside {[3:5]};  // Multiple reset events
  }) begin
    `uvm_error(get_type_name(), "Failed to randomize reset sequence")
  end
  
  `uvm_info(get_type_name(), $sformatf("Testing with %0d reset events", reset_seq.num_reset_events), UVM_LOW)
  
  if (test_config.num_masters > 0) begin
    reset_seq.start(axi4_env_h.axi4_virtual_seqr_h.axi4_master_write_seqr_h_all[0]);
  end else begin
    reset_seq.start(axi4_env_h.axi4_virtual_seqr_h.axi4_master_write_seqr_h);
  end
  
  // Wait for completion
  #500ns;
  
  phase.drop_objection(this);
  
endtask : run_phase

//--------------------------------------------------------------------------------------------
// Class: axi4_exception_clk_reset_combined_test
// Description:
// This test combines clock frequency changes and reset termination.
// - Mixed exceptions: Clock changes, resets, or both simultaneous
// - Number of events: 3-15 (random)
// - Tests system resilience under combined stress
// - Verifies proper recovery and protocol compliance
// - Supports all bus matrix modes (NONE/1x1, BASE/4x4, ENHANCED/10x10)
//--------------------------------------------------------------------------------------------
class axi4_exception_clk_reset_combined_test extends axi4_error_inject_base_test;
  `uvm_component_utils(axi4_exception_clk_reset_combined_test)

  extern function new(string name = "axi4_exception_clk_reset_combined_test", uvm_component parent = null);
  extern function void build_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);

endclass : axi4_exception_clk_reset_combined_test

function axi4_exception_clk_reset_combined_test::new(string name = "axi4_exception_clk_reset_combined_test", uvm_component parent = null);
  super.new(name, parent);
endfunction : new

function void axi4_exception_clk_reset_combined_test::build_phase(uvm_phase phase);
  super.build_phase(phase);
  
  // Configure test for combined clock and reset exceptions
  uvm_config_db#(bit)::set(this, "*", "enable_exceptions", 1);
  uvm_config_db#(bit)::set(this, "*", "clk_freq_exception", 1);
  uvm_config_db#(bit)::set(this, "*", "reset_terminate", 1);
  uvm_config_db#(bit)::set(this, "*", "combined_exceptions", 1);
  
  `uvm_info(get_type_name(), "Build phase completed for Combined Clock/Reset test", UVM_LOW)
endfunction : build_phase

task axi4_exception_clk_reset_combined_test::run_phase(uvm_phase phase);
  axi4_virtual_exception_clk_reset_seq combined_seq;
  
  phase.raise_objection(this);
  
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  `uvm_info(get_type_name(), "Starting Combined Clock/Reset Exception Test", UVM_LOW)
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  `uvm_info(get_type_name(), "Test Description:", UVM_LOW)
  `uvm_info(get_type_name(), "  - Mixed clock and reset exceptions", UVM_LOW)
  `uvm_info(get_type_name(), "  - Simultaneous exception events", UVM_LOW)
  `uvm_info(get_type_name(), "  - Tests combined stress scenarios", UVM_LOW)
  `uvm_info(get_type_name(), $sformatf("  - Bus Matrix Mode: %s with %0dx%0d configuration", 
            test_config.bus_matrix_mode.name(), test_config.num_masters, test_config.num_slaves), UVM_LOW)
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  
  // Run the combined exception sequence
  combined_seq = axi4_virtual_exception_clk_reset_seq::type_id::create("combined_seq");
  combined_seq.start(axi4_env_h.axi4_virtual_seqr_h);
  
  // Wait for completion
  #2000ns;
  
  phase.drop_objection(this);
  
endtask : run_phase

//--------------------------------------------------------------------------------------------
// Class: axi4_exception_continuous_clk_change_test
// Description:
// This test continuously changes clock frequency throughout simulation.
// - Continuous frequency variation: 5-30% probability per interval
// - Test duration: 5-20 us
// - Random frequency factors: 0.5x to 3.0x
// - Background traffic during changes
// - Supports all bus matrix modes (NONE/1x1, BASE/4x4, ENHANCED/10x10)
//--------------------------------------------------------------------------------------------
class axi4_exception_continuous_clk_change_test extends axi4_error_inject_base_test;
  `uvm_component_utils(axi4_exception_continuous_clk_change_test)

  extern function new(string name = "axi4_exception_continuous_clk_change_test", uvm_component parent = null);
  extern function void build_phase(uvm_phase phase);
  extern virtual function void setup_axi4_env_cfg();
  extern task run_phase(uvm_phase phase);

endclass : axi4_exception_continuous_clk_change_test

function axi4_exception_continuous_clk_change_test::new(string name = "axi4_exception_continuous_clk_change_test", uvm_component parent = null);
  super.new(name, parent);
endfunction : new

function void axi4_exception_continuous_clk_change_test::build_phase(uvm_phase phase);
  super.build_phase(phase);
  
  // Configure test for continuous clock frequency changes
  uvm_config_db#(bit)::set(this, "*", "enable_exceptions", 1);
  uvm_config_db#(bit)::set(this, "*", "continuous_clk_change", 1);
  uvm_config_db#(int)::set(this, "*", "clk_change_probability", 15);  // 15% chance
  
  `uvm_info(get_type_name(), "Build phase completed for Continuous Clock Change test", UVM_LOW)
endfunction : build_phase

function void axi4_exception_continuous_clk_change_test::setup_axi4_env_cfg();
  // Call parent implementation first
  super.setup_axi4_env_cfg();
  
  // Enable frequency checker for this test
  axi4_env_cfg_h.has_freq_checker = 1;
  
  // Configure expected frequency changes for the checker
  // The test performs about 20 random frequency changes with 15% probability
  uvm_config_db#(int)::set(this, "*", "expected_freq_changes", 20);
  
  `uvm_info(get_type_name(), "Enabled frequency checker for continuous clock change test", UVM_MEDIUM)
endfunction : setup_axi4_env_cfg

task axi4_exception_continuous_clk_change_test::run_phase(uvm_phase phase);
  axi4_master_exception_clk_freq_seq clk_seq;
  axi4_master_write_seq write_seq;
  int freq_idx;
  int active_masters;
  int total_freq_changes = 0;
  
  phase.raise_objection(this);
  
  // Determine active masters based on bus matrix mode
  case(test_config.bus_matrix_mode)
    axi4_bus_matrix_ref::NONE: active_masters = 1;
    axi4_bus_matrix_ref::BASE_BUS_MATRIX: active_masters = 4;
    axi4_bus_matrix_ref::BUS_ENHANCED_MATRIX: active_masters = test_config.num_masters;
  endcase
  
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  `uvm_info(get_type_name(), "Starting Continuous Clock Change Test", UVM_LOW)
  `uvm_info(get_type_name(), $sformatf("  Active Masters: %0d", active_masters), UVM_LOW)
  `uvm_info(get_type_name(), "===============================================", UVM_LOW)
  
  // Configure expected frequency changes for the checker
  if(axi4_env_h.axi4_freq_checker_h != null) begin
    // Don't set strict expectations, just monitor
    axi4_env_h.axi4_freq_checker_h.expected_freq_changes = 0;  // 0 means no strict checking
  end
  
  // Run continuous clock changes with background traffic on multiple interfaces
  fork
    // Background traffic on all active masters
    begin
      for(int m = 0; m < active_masters; m++) begin
        automatic int master_id = m;
        fork
          begin
            repeat(50) begin
              write_seq = axi4_master_write_seq::type_id::create($sformatf("write_seq_m%0d", master_id));
              if(!write_seq.randomize()) begin
                `uvm_error(get_type_name(), $sformatf("Write sequence randomization failed for master %0d", master_id))
              end
              if (test_config.num_masters > master_id) begin
                write_seq.start(axi4_env_h.axi4_virtual_seqr_h.axi4_master_write_seqr_h_all[master_id]);
              end
              #40ns;
            end
          end
        join_none
      end
    end
    
    // Continuous clock changes on different interfaces
    begin
      repeat(20) begin
        if ($urandom_range(0, 100) < 15) begin  // 15% probability
          int target_master = $urandom_range(0, active_masters-1);
          freq_idx = $urandom_range(0, 6);  // 0-6 for scale factor index
          
          `uvm_info(get_type_name(), $sformatf("Changing frequency for master %0d to scale index %0d", 
                    target_master, freq_idx), UVM_MEDIUM)
          
          clk_seq = axi4_master_exception_clk_freq_seq::type_id::create($sformatf("clk_seq_m%0d", target_master));
          if(!clk_seq.randomize() with {
            num_freq_changes == 1;
            freq_scale_idx[0] == local::freq_idx;
            freq_hold_cycles[0] inside {[10:50]};
          }) begin
            `uvm_error(get_type_name(), "Clock sequence randomization failed")
          end
          
          if (test_config.num_masters > target_master) begin
            clk_seq.start(axi4_env_h.axi4_virtual_seqr_h.axi4_master_write_seqr_h_all[target_master]);
          end
          
          total_freq_changes++;
        end
        #100ns;
      end
    end
  join
  
  `uvm_info(get_type_name(), $sformatf("Total frequency changes: %0d", total_freq_changes), UVM_LOW)
  
  phase.drop_objection(this);
  
endtask : run_phase

`endif