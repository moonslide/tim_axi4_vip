class c_43_9;
    bit[63:0] awaddr = 64'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../slave/axi4_slave_driver_proxy.sv:222)
    {
       (awaddr != 0);
    }
endclass

program p_43_9;
    c_43_9 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x00x1z0000z0xxz0010xxzz0zz0xx0x0zxxxzxzxxxxzxxzzzxzxxzzzxzzxzxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
