`ifndef AXI4_QOS_STARVATION_PREVENTION_TEST_INCLUDED_
`define AXI4_QOS_STARVATION_PREVENTION_TEST_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: axi4_qos_starvation_prevention_test
// 
// TEST SCENARIO DESCRIPTION:
// ==========================
// This test validates that the QoS arbitration system prevents indefinite starvation
// of low priority transactions when high priority traffic is continuously present.
// It verifies that fairness mechanisms ensure all transactions eventually get serviced
// within reasonable time bounds.
//
// DETAILED TEST SCENARIOS:
// 1. Continuous High Priority vs Low Priority Test:
//    - Master 0: Generates continuous high priority transactions (QoS 0xF)
//    - Master 1: Generates low priority transactions (QoS 0x0)
//    - Validates that low priority transactions are not indefinitely blocked
//    - Measures maximum response time for low priority transactions
//
// 2. Mixed Priority Starvation Test:
//    - Master 0: High priority (QoS 0xF) - 60% of traffic
//    - Master 1: Medium priority (QoS 0x8) - 30% of traffic
//    - Master 2: Low priority (QoS 0x2) - 10% of traffic
//    - Tests proportional fairness with aging mechanisms
//    - Ensures lowest priority gets minimum guaranteed service
//
// 3. Temporal Priority Escalation Test:
//    - Low priority transactions that age beyond threshold get priority boost
//    - Tests aging algorithms that prevent starvation
//    - Validates that aged transactions receive elevated service
//    - Measures effectiveness of temporal priority escalation
//
// 4. Burst-Induced Starvation Test:
//    - High priority master generates large bursts (AWLEN=15) continuously
//    - Low priority master generates single-beat transactions
//    - Tests fairness when high priority consumes significant resources
//    - Validates that resource consumption doesn't cause indefinite starvation
//
// 5. Multi-Slave Starvation Prevention Test:
//    - High priority traffic targets Slave 0
//    - Low priority traffic targets Slave 1
//    - Mixed priority traffic targets Slave 2
//    - Validates starvation prevention across different slave interfaces
//    - Ensures per-slave fairness mechanisms work correctly
//
// STARVATION SCENARIOS:
// - Continuous high priority traffic generation
// - Resource-intensive high priority transactions (large bursts)
// - Multiple high priority masters vs single low priority master
// - Worst-case timing patterns designed to expose starvation
//
// EXPECTED BEHAVIORS:
// - Low priority transactions should complete within bounded time
// - Maximum starvation time should not exceed system-defined thresholds
// - High priority transactions should maintain their precedence
// - Aging mechanisms should escalate long-waiting transactions
// - System should maintain fairness while respecting priority ordering
//
// STARVATION PREVENTION MECHANISMS:
// - Temporal aging algorithms that boost priority over time
// - Minimum service guarantees for low priority traffic
// - Round-robin fairness within same priority levels
// - Bounded waiting time limits with escalation policies
// - Resource reservation for low priority transactions
//
// METRICS:
// - Maximum response time for each priority level
// - Starvation duration measurements
// - Fairness index calculations
// - Priority escalation event tracking
// - Service ratio analysis across priority levels
//
// COVERAGE GOALS:
// - All priority level combinations and interactions
// - Starvation prevention mechanism activation
// - Temporal aging and priority escalation events
// - Bounded waiting time validation
// - Multi-slave fairness verification
//--------------------------------------------------------------------------------------------
class axi4_qos_starvation_prevention_test extends axi4_base_test;
  `uvm_component_utils(axi4_qos_starvation_prevention_test)
  
  // Virtual sequence handle
  axi4_virtual_qos_starvation_prevention_seq axi4_virtual_qos_starvation_prevention_seq_h;
  
  //-------------------------------------------------------
  // Externally defined Tasks and Functions
  //-------------------------------------------------------
  extern function new(string name = "axi4_qos_starvation_prevention_test", uvm_component parent = null);
  extern virtual function void build_phase(uvm_phase phase);
  extern virtual task run_phase(uvm_phase phase);
  
endclass : axi4_qos_starvation_prevention_test

//--------------------------------------------------------------------------------------------
// Construct: new
//--------------------------------------------------------------------------------------------
function axi4_qos_starvation_prevention_test::new(string name = "axi4_qos_starvation_prevention_test", uvm_component parent = null);
  super.new(name, parent);
endfunction : new

//--------------------------------------------------------------------------------------------
// Function: build_phase
// Creates test configuration and components
//--------------------------------------------------------------------------------------------
function void axi4_qos_starvation_prevention_test::build_phase(uvm_phase phase);
  // Set configuration before calling super.build_phase()
  `uvm_info(get_type_name(), "Configuring QoS starvation prevention test", UVM_MEDIUM)
  
  super.build_phase(phase);
  
  // Enable QoS mode for all agents in QoS tests
  for (int i = 0; i < axi4_env_cfg_h.no_of_masters; i++) begin
    axi4_env_cfg_h.axi4_master_agent_cfg_h[i].qos_mode_type = WRITE_READ_QOS_MODE_ENABLE;
  end
  for (int i = 0; i < axi4_env_cfg_h.no_of_slaves; i++) begin
    axi4_env_cfg_h.axi4_slave_agent_cfg_h[i].qos_mode_type = WRITE_READ_QOS_MODE_ENABLE;
  end
  `uvm_info(get_type_name(), "Enabled WRITE_READ_QOS_MODE for all agents", UVM_LOW)
  
  // Set reasonable timeout for starvation prevention test
  uvm_top.set_timeout(30ms, 0); // 30ms timeout for starvation test
  
  // Set enhanced bus matrix mode for QoS testing  
  test_config.bus_matrix_mode = axi4_bus_matrix_ref::BUS_ENHANCED_MATRIX;
  
  // Update config_db with the correct bus matrix mode
  uvm_config_db#(axi4_bus_matrix_ref::bus_matrix_mode_e)::set(this, "*", "bus_matrix_mode", test_config.bus_matrix_mode);
  
  `uvm_info(get_type_name(), "QoS starvation prevention test configuration completed", UVM_MEDIUM)
  
endfunction : build_phase

//--------------------------------------------------------------------------------------------
// Task: run_phase
// Executes the QoS starvation prevention test
//--------------------------------------------------------------------------------------------
task axi4_qos_starvation_prevention_test::run_phase(uvm_phase phase);
  
  phase.raise_objection(this, "axi4_qos_starvation_prevention_test");
  
  `uvm_info(get_type_name(), "Starting AXI4 QoS Starvation Prevention Test", UVM_LOW)
  `uvm_info(get_type_name(), "Test objective: Verify low priority traffic is not starved by high priority traffic", UVM_LOW)
  
  // Create and start the virtual sequence
  axi4_virtual_qos_starvation_prevention_seq_h = axi4_virtual_qos_starvation_prevention_seq::type_id::create("axi4_virtual_qos_starvation_prevention_seq_h");
  
  // Configure the virtual sequence  
  axi4_virtual_qos_starvation_prevention_seq_h.start(axi4_env_h.axi4_virtual_seqr_h);
  
  // Wait for all transactions to complete, including low priority ones
  #8000;
  
  `uvm_info(get_type_name(), "AXI4 QoS Starvation Prevention Test completed", UVM_LOW)
  `uvm_info(get_type_name(), "Test success criteria:", UVM_LOW)
  `uvm_info(get_type_name(), "1. All low priority transactions eventually completed", UVM_LOW)
  `uvm_info(get_type_name(), "2. High priority transactions maintained precedence", UVM_LOW)
  `uvm_info(get_type_name(), "3. No indefinite starvation occurred", UVM_LOW)
  `uvm_info(get_type_name(), "4. Fair arbitration was demonstrated", UVM_LOW)
  `uvm_info(get_type_name(), "5. Maximum response time bounds were respected", UVM_LOW)
  
  phase.drop_objection(this, "axi4_qos_starvation_prevention_test");
  
endtask : run_phase

`endif