`ifndef AXI4_QOS_EQUAL_PRIORITY_FAIRNESS_TEST_INCLUDED_
`define AXI4_QOS_EQUAL_PRIORITY_FAIRNESS_TEST_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: axi4_qos_equal_priority_fairness_test
// 
// TEST SCENARIO DESCRIPTION:
// ==========================
// This test validates fair arbitration and bandwidth allocation when multiple masters 
// generate transactions with identical QoS values. It ensures that no master is starved
// and that bandwidth is distributed equitably among competing masters.
//
// DETAILED TEST SCENARIOS:
// 1. Equal QoS Fair Arbitration Test:
//    - 4 masters simultaneously generate transactions with identical QoS (0x8)
//    - Each master generates 50 transactions targeting the same slave
//    - Validates round-robin or weighted fair queuing arbitration
//    - Measures bandwidth allocation per master for fairness analysis
//
// 2. Sustained Equal Priority Load Test:
//    - Continuous transaction generation with equal QoS across all masters
//    - Tests system behavior under sustained equal-priority contention
//    - Validates that no master experiences significant delays relative to others
//    - Measures average latency and throughput per master
//
// 3. Mixed Transaction Types Fairness Test:
//    - Masters generate both read and write transactions with equal QoS
//    - Even masters: Write-focused workload (70% writes, 30% reads)
//    - Odd masters: Read-focused workload (30% writes, 70% reads)
//    - Validates fairness across different transaction types
//
// 4. Burst Length Fairness Test:
//    - Masters generate transactions with varying burst lengths but equal QoS
//    - Master 0: Short bursts (1-2 beats)
//    - Master 1: Medium bursts (4-8 beats)  
//    - Master 2: Long bursts (8-16 beats)
//    - Master 3: Mixed burst lengths
//    - Ensures fairness regardless of burst length differences
//
// EXPECTED BEHAVIORS:
// - Each master should receive approximately equal bandwidth allocation
// - No master should be completely starved for extended periods
// - Arbitration should be deterministic and predictable
// - Total system throughput should be maximized while maintaining fairness
// - Latency variation between masters should be minimal
//
// FAIRNESS METRICS:
// - Bandwidth allocation deviation should be < 10% between masters
// - Maximum starvation time should be bounded and reasonable
// - Transaction completion rate should be similar across masters
// - Jitter in service intervals should be minimized
//
// COVERAGE GOALS:
// - Equal QoS arbitration algorithms (round-robin, weighted fair queuing)
// - Sustained contention scenarios
// - Mixed workload fairness validation
// - Bandwidth allocation measurement and analysis
// 
// Uses enhanced 4x4 bus matrix configuration (scaled from 10x10 specification)
//--------------------------------------------------------------------------------------------
class axi4_qos_equal_priority_fairness_test extends axi4_base_test;
  
  `uvm_component_utils(axi4_qos_equal_priority_fairness_test)
  
  // Virtual sequence handle
  axi4_virtual_qos_equal_priority_fairness_seq qos_fairness_vseq;
  
  //-------------------------------------------------------
  // Externally defined tasks and functions
  //-------------------------------------------------------
  extern function new(string name = "axi4_qos_equal_priority_fairness_test", uvm_component parent = null);
  extern virtual function void build_phase(uvm_phase phase);
  extern virtual task run_phase(uvm_phase phase);
  
endclass : axi4_qos_equal_priority_fairness_test

//-----------------------------------------------------------------------------
// Constructor: new
//-----------------------------------------------------------------------------
function axi4_qos_equal_priority_fairness_test::new(string name = "axi4_qos_equal_priority_fairness_test", uvm_component parent = null);
  super.new(name, parent);
endfunction : new

//-----------------------------------------------------------------------------
// Function: build_phase
// Configure the test for 10x10 enhanced bus matrix
//-----------------------------------------------------------------------------
function void axi4_qos_equal_priority_fairness_test::build_phase(uvm_phase phase);
  // Set configuration before calling super.build_phase()
  `uvm_info(get_type_name(), "Configuring QoS equal priority fairness test", UVM_LOW)
  
  // Create and configure test_config BEFORE calling super.build_phase()
  test_config = axi4_test_config::type_id::create("test_config");
  test_config.configure_for_test(get_type_name());
  
  // Ensure we're using 10x10 configuration for this test BEFORE calling super.build_phase()
  if (test_config.num_masters < 10 || test_config.num_slaves < 10) begin
    `uvm_warning(get_type_name(), "QoS test designed for 10x10 bus matrix. Adjusting configuration.")
    test_config.num_masters = 10;
    test_config.num_slaves = 10;
  end
  
  // Set enhanced bus matrix mode for QoS testing BEFORE calling super.build_phase()
  test_config.bus_matrix_mode = axi4_bus_matrix_ref::BUS_ENHANCED_MATRIX;
  
  `uvm_info(get_type_name(), $sformatf("QoS test config override: bus_matrix_mode=%s, masters=%0d, slaves=%0d", 
                                       test_config.bus_matrix_mode.name(), test_config.num_masters, test_config.num_slaves), UVM_LOW)
  
  // Store in config_db for use by environment and other components
  uvm_config_db#(axi4_test_config)::set(this, "*", "test_config", test_config);
  uvm_config_db#(axi4_bus_matrix_ref::bus_matrix_mode_e)::set(this, "*", "bus_matrix_mode", test_config.bus_matrix_mode);
  
  super.build_phase(phase);
  
  // Enable QoS mode for all agents in QoS tests
  for (int i = 0; i < axi4_env_cfg_h.no_of_masters; i++) begin
    axi4_env_cfg_h.axi4_master_agent_cfg_h[i].qos_mode_type = WRITE_READ_QOS_MODE_ENABLE;
  end
  for (int i = 0; i < axi4_env_cfg_h.no_of_slaves; i++) begin
    axi4_env_cfg_h.axi4_slave_agent_cfg_h[i].qos_mode_type = WRITE_READ_QOS_MODE_ENABLE;
  end
  `uvm_info(get_type_name(), "Enabled WRITE_READ_QOS_MODE for all agents", UVM_LOW)
  
  // Force proper slave configuration for QoS tests regardless of auto-configuration
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[0].min_address = 64'h0000_0008_0000_0000;
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[0].max_address = 64'h0000_0008_3FFF_FFFF;
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[1].min_address = 64'h0000_0008_4000_0000;
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[1].max_address = 64'h0000_0008_7FFF_FFFF;
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[2].min_address = 64'h0000_0008_8000_0000;
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[2].max_address = 64'h0000_0008_BFFF_FFFF;
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[3].min_address = 64'h0000_0008_C000_0000;
  axi4_env_cfg_h.axi4_slave_agent_cfg_h[3].max_address = 64'h0000_0008_FFFF_FFFF;
  
  // Set higher timeout for this longer test
  uvm_config_db#(time)::set(this, "*", "timeout", 500ms);
  
  // Set timeout for equal priority fairness test with random masters
  uvm_top.set_timeout(20ms, 0); // 20ms timeout for random master configs
  
endfunction : build_phase

//-----------------------------------------------------------------------------
// Task: run_phase
// Run the QoS equal priority fairness virtual sequence
//-----------------------------------------------------------------------------
task axi4_qos_equal_priority_fairness_test::run_phase(uvm_phase phase);
  
  `uvm_info(get_type_name(), "Starting QoS equal priority fairness test", UVM_MEDIUM)
  
  // Create the virtual sequence
  qos_fairness_vseq = axi4_virtual_qos_equal_priority_fairness_seq::type_id::create("qos_fairness_vseq");
  
  phase.raise_objection(this);
  
  // Start the virtual sequence
  qos_fairness_vseq.start(axi4_env_h.axi4_virtual_seqr_h);
  
  // Add extra time for scoreboard checking and bandwidth measurement
  #10000;
  
  phase.drop_objection(this);
  
  `uvm_info(get_type_name(), "QoS equal priority fairness test completed", UVM_MEDIUM)
  `uvm_info(get_type_name(), "Check simulation logs for bandwidth allocation statistics", UVM_MEDIUM)
  
endtask : run_phase

`endif