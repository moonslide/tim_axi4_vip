`ifndef AXI4_SLAVE_MEMORY_INCLUDED_
`define AXI4_SLAVE_MEMORY_INCLUDED_

import axi4_config_pkg::*;

//--------------------------------------------------------------------------------------------
// Class: axi4_slave_agent
// This agent has sequencer, driver_proxy, monitor_proxy for axi4  
//--------------------------------------------------------------------------------------------
class axi4_slave_memory extends uvm_object;
  `uvm_object_utils(axi4_slave_memory)

  import axi4_config_pkg::*;

  // uvm_mem model for this slave
  uvm_mem mem;
  // Base address used for index calculations
  bit [ADDRESS_WIDTH-1:0] base_addr;

  //Variable : slave_memory
  //Declaration of slave_memory to store the data from master
  protected bit [7:0] slave_memory [longint];

  //Variable : fifo_memory
  //Declaration of fifo_memory to store the data from master of type fixed
  protected bit [7:0] fifo_memory [$];

  extern function new(string name = "axi4_slave_memory");  
  extern virtual function void mem_write(input bit [ADDRESS_WIDTH-1:0]slave_address,
                                         bit [DATA_WIDTH-1:0] data);
  extern virtual function void mem_read (input bit [ADDRESS_WIDTH-1:0]slave_address,
                                         output bit [DATA_WIDTH-1:0] data);
  extern virtual function void fifo_write(input bit [DATA_WIDTH-1:0]data);
  extern virtual function void fifo_read (output bit [DATA_WIDTH-1:0]data);
  extern virtual function bit is_slave_addr_exists(input bit [ADDRESS_WIDTH-1 :0]slave_address);
  extern static function string get_slave_for_address(bit [ADDRESS_WIDTH-1:0] addr);
  extern static function bit    master_has_access(string mname, string sname);

endclass : axi4_slave_memory

//--------------------------------------------------------------------------------------------
// Construct: new
//
// Parameters:
//  name - axi4_slave_agent_config
//--------------------------------------------------------------------------------------------
function axi4_slave_memory::new(string name = "axi4_slave_memory");
  super.new(name);
  // Determine base address for this memory based on name
  foreach(slave_addr_table[i]) begin
    if(slave_addr_table[i].slave_name == name) begin
      base_addr = slave_addr_table[i].base_addr;
      mem = new(name,
                slave_addr_table[i].size/STROBE_WIDTH,
                DATA_WIDTH,
                "RW");
    end
  end
endfunction : new


//--------------------------------------------------------------------------------------------
//Task : mem_write
//Used to store the slave data into the slave memory
//Parameter :
//slave_address - bit [ADDRESS_WIDTH-1 :0]
//data          - bit [DATA_WIDTH-1:0]
//--------------------------------------------------------------------------------------------
function void axi4_slave_memory::mem_write(input bit [ADDRESS_WIDTH-1 :0]slave_address,
                                           bit [DATA_WIDTH-1:0] data);
  slave_memory[slave_address] = data;
  if(mem != null) begin
    int unsigned idx = (slave_address - base_addr)/STROBE_WIDTH;
    mem.poke(idx, data);
  end
endfunction : mem_write

//--------------------------------------------------------------------------------------------
//Task : mem_read
//Used to store the slave data into the slave memory
//Parameter :
//slave_address - bit [ADDRESS_WIDTH-1 :0]
//data          - bit [DATA_WIDTH-1:0]
//--------------------------------------------------------------------------------------------
function void axi4_slave_memory::mem_read(input bit [ADDRESS_WIDTH-1 :0]slave_address,
                                          output bit [DATA_WIDTH-1:0] data);
  if(mem != null) begin
    int unsigned idx = (slave_address - base_addr)/STROBE_WIDTH;
    mem.peek(idx, data);
  end
  else begin
    data = slave_memory[slave_address];
  end
endfunction : mem_read

//--------------------------------------------------------------------------------------------
//Task : fifo_write
//Used to store the slave data into the slave memory
//Parameter :
//data          - bit [DATA_WIDTH-1:0]
//--------------------------------------------------------------------------------------------
function void axi4_slave_memory::fifo_write(input bit [DATA_WIDTH-1:0]data);
  fifo_memory.push_front(data);
endfunction : fifo_write

//--------------------------------------------------------------------------------------------
//Task : fifo_read
//Used to store the slave data into the slave memory
//Parameter :
//data          - bit [DATA_WIDTH-1:0]
//--------------------------------------------------------------------------------------------
function void axi4_slave_memory::fifo_read(output bit [DATA_WIDTH-1:0]data);
  data = fifo_memory.pop_back();
endfunction : fifo_read

//--------------------------------------------------------------------------------------------
//Task : is_slave_addr_exists
//Used to check the address exists are not in the memory
//slave_address - bit [ADDRESS_WIDTH-1 :0]
//--------------------------------------------------------------------------------------------
function bit axi4_slave_memory::is_slave_addr_exists(input bit [ADDRESS_WIDTH-1 :0]slave_address);
  if(mem != null) begin
    int unsigned idx = (slave_address - base_addr)/STROBE_WIDTH;
    bit [DATA_WIDTH-1:0] tmp;
    mem.peek(idx, tmp);
    is_slave_addr_exists = 1;
  end
  else begin
    is_slave_addr_exists = slave_memory.exists(slave_address);
  end
endfunction: is_slave_addr_exists

// Return slave name for an address
static function string axi4_slave_memory::get_slave_for_address(bit [ADDRESS_WIDTH-1:0] addr);
  foreach(slave_addr_table[i]) begin
    if(addr >= slave_addr_table[i].base_addr && addr < slave_addr_table[i].base_addr + slave_addr_table[i].size)
      return slave_addr_table[i].slave_name;
  end
  return "";
endfunction

// Check if a master is allowed to access a slave
static function bit axi4_slave_memory::master_has_access(string mname, string sname);
  foreach(master_access_table[i]) begin
    if(master_access_table[i].master_name == mname) begin
      foreach(master_access_table[i].allowed_slaves[j])
        if(master_access_table[i].allowed_slaves[j] == sname)
          return 1;
    end
  end
  return 0;
endfunction


`endif
