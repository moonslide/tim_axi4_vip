class c_41_9;
    bit[63:0] awaddr = 64'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../slave/axi4_slave_driver_proxy.sv:222)
    {
       (awaddr != 0);
    }
endclass

program p_41_9;
    c_41_9 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zx0z0xz00x1000zzzz1z1z111xzxx111zxxzxxxzzzxxzzzxxzxzxxxzxzzzxxxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
