class c_52_9;
    bit[63:0] awaddr = 64'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../slave/axi4_slave_driver_proxy.sv:222)
    {
       (awaddr != 0);
    }
endclass

program p_52_9;
    c_52_9 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "x0xzx1011xxzxx01xx0xxz00101x110xxzxzzzxzxxxxxxzzzxxzxzzzzzxxxxzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
