class c_35_9;
    bit[63:0] awaddr = 64'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../slave/axi4_slave_driver_proxy.sv:222)
    {
       (awaddr != 0);
    }
endclass

program p_35_9;
    c_35_9 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z11zx11x101zx1x0x111zxz1x1x1xzzxxzxxxzxxxzxzxxzxzxzzzxzxzxzzxxzx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
