`ifndef AXI4_BUS_MATRIX_PKG_INCLUDED_
`define AXI4_BUS_MATRIX_PKG_INCLUDED_
package axi4_bus_matrix_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import axi4_globals_pkg::*;
  import axi4_slave_pkg::*;
  `include "axi4_bus_matrix_ref.sv"
endpackage : axi4_bus_matrix_pkg
`endif
