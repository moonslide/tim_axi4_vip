class c_5_9;
    bit[63:0] awaddr = 64'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../slave/axi4_slave_driver_proxy.sv:222)
    {
       (awaddr != 0);
    }
endclass

program p_5_9;
    c_5_9 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "1zxz11zxz000011xxxxzxz1zz1zxzz00zxzzxxxxzzzxxxzxzxzxzzxxxxzzzzzz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
