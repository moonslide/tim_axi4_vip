class c_26_9;
    bit[63:0] awaddr = 64'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../slave/axi4_slave_driver_proxy.sv:222)
    {
       (awaddr != 0);
    }
endclass

program p_26_9;
    c_26_9 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "zzz0zzzx1z0zzx0x00x1xxxz0110xx01zxxxzzxxzxxxxxxxzxxzzxzzxzxzzzxx";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
