class c_50_9;
    bit[63:0] awaddr = 64'h0;

    constraint WITH_CONSTRAINT_this    // (constraint_mode = ON) (../slave/axi4_slave_driver_proxy.sv:222)
    {
       (awaddr != 0);
    }
endclass

program p_50_9;
    c_50_9 obj;
    string randState;

    initial
        begin
            obj = new;
            randState = "z10zx1x111x000011xzxx0zzz01x0010xzxzxzxzzxzzzxxxxxxxzxxxzzzxxzxz";
            obj.set_randstate(randState);
            obj.randomize();
        end
endprogram
