`ifndef AXI4_MASTER_QOS_WRITE_ONLY_SEQ_INCLUDED_
`define AXI4_MASTER_QOS_WRITE_ONLY_SEQ_INCLUDED_

//--------------------------------------------------------------------------------------------
// Class: axi4_master_qos_write_only_seq
// Dedicated write-only sequence for QoS equal priority fairness test
// This sequence ONLY generates WRITE transactions
//--------------------------------------------------------------------------------------------
class axi4_master_qos_write_only_seq extends axi4_master_base_seq;

  `uvm_object_utils(axi4_master_qos_write_only_seq)
  
  // Transaction handle
  axi4_master_tx req;
  
  // Master and slave IDs for this sequence
  int master_id;
  int slave_id;
  
  // Test parameters
  bit [3:0] qos_value = 4'h8; // All masters use same QoS
  int num_transactions = 1;   // Minimal transactions for basic functionality testing
  int inter_transaction_delay = 100; // Reduced delay for faster completion
  
  // Transaction ID counter to ensure unique IDs per sequence instance
  int unsigned transaction_id_counter = 0;
  
  //-------------------------------------------------------
  // Externally defined tasks and functions
  //-------------------------------------------------------
  extern function new(string name = "axi4_master_qos_write_only_seq");
  extern virtual task body();
  extern function bit [ADDRESS_WIDTH-1:0] calculate_slave_address(int slave_id);
  
endclass : axi4_master_qos_write_only_seq

//-----------------------------------------------------------------------------
// Constructor: new
//-----------------------------------------------------------------------------
function axi4_master_qos_write_only_seq::new(string name = "axi4_master_qos_write_only_seq");
  super.new(name);
endfunction : new

//-----------------------------------------------------------------------------
// Task: body
// Main sequence body - generates WRITE transactions ONLY
//-----------------------------------------------------------------------------
task axi4_master_qos_write_only_seq::body();
  bit [15:0] calculated_id;
  super.body();
  
  // Get master and slave IDs from configuration
  if (!uvm_config_db#(int)::get(null, get_full_name(), "master_id", master_id)) begin
    master_id = 0; // Default to even master ID for write
  end
  
  if (!uvm_config_db#(int)::get(null, get_full_name(), "slave_id", slave_id)) begin
    slave_id = 2; // Default to slave 2
  end
  
  // Minimal stagger delay 
  #(master_id * 100ns);
  
  // Get test parameters from config if available
  void'(uvm_config_db#(bit [3:0])::get(null, get_full_name(), "qos_value", qos_value));
  void'(uvm_config_db#(int)::get(null, get_full_name(), "num_transactions", num_transactions));
  
  `uvm_info(get_type_name(), $sformatf("Starting WRITE-ONLY QoS sequence - Master %0d to Slave %0d with QoS=0x%0h", 
                                       master_id, slave_id, qos_value), UVM_MEDIUM)
  
  // Generate WRITE transactions ONLY
  for (int i = 0; i < num_transactions; i++) begin
    // Create and send write transaction using proper UVM sequence protocol
    req = axi4_master_tx::type_id::create("req");
    
    // Calculate unique ID within 16-value constraint
    // Use master_id as base and add transaction counter modulo (16-master_id) to avoid overlap
    calculated_id = master_id + (transaction_id_counter % (16 - master_id));
    if (calculated_id >= 16) calculated_id = master_id; // Wrap around if needed
    if (calculated_id == 0) calculated_id = 1; // Avoid ID 0
    
    start_item(req);
    if(!req.randomize() with {
      req.tx_type == WRITE;
      req.awaddr == calculate_slave_address(slave_id) + (i * 'h1000) + (master_id * 'h100);
      req.awid == `GET_AWID_ENUM(calculated_id);
      req.awlen == 0;  // Force single-beat transactions only
      req.awsize == WRITE_8_BYTES;
      req.awburst == WRITE_INCR;
      req.awqos == qos_value;
      // Ensure read address is a valid slave address for write transactions to avoid DECERR
      req.araddr == 64'h0000_0008_0000_0000;
    }) begin
      `uvm_error(get_type_name(), "Failed to randomize write transaction")
    end
    transaction_id_counter++;
    
    finish_item(req);
    
    // Minimal inter-transaction delay 
    #(inter_transaction_delay * 10ns);
  end
  
  `uvm_info(get_type_name(), $sformatf("WRITE-ONLY QoS sequence completed - sent %0d write transactions", num_transactions), UVM_MEDIUM)
  
endtask : body

//-----------------------------------------------------------------------------
// Function: calculate_slave_address
// Calculate base address for slave based on slave ID
//-----------------------------------------------------------------------------
function bit [ADDRESS_WIDTH-1:0] axi4_master_qos_write_only_seq::calculate_slave_address(int slave_id);
  // Enhanced bus matrix address mapping - must match axi4_bus_matrix_ref.sv configuration
  case(slave_id)
    0: return 64'h0000_0008_0000_0000; // S0: DDR Secure Kernel
    1: return 64'h0000_0008_4000_0000; // S1: DDR Non-Secure User
    2: return 64'h0000_0008_8000_0000; // S2: DDR Shared Buffer
    3: return 64'h0000_0008_C000_0000; // S3: Illegal Address Hole (will return DECERR)
    4: return 64'h0000_0009_0000_0000; // S4: XOM Instruction-Only (read-only, will return SLVERR on write)
    5: return 64'h0000_000A_0000_0000; // S5: RO Peripheral (read-only, will return SLVERR on write)
    6: return 64'h0000_000A_0001_0000; // S6: Privileged-Only
    7: return 64'h0000_000A_0002_0000; // S7: Secure-Only
    8: return 64'h0000_000A_0003_0000; // S8: Scratchpad
    9: return 64'h0000_000A_0004_0000; // S9: Attribute Monitor
    default: return 64'h0000_0008_8000_0000; // Default to S2: DDR Shared Buffer
  endcase
endfunction : calculate_slave_address

`endif